cw7800

.SUBCKT LM7805C 19 8 21
QAP 4 3 19 QPMOD
Q1N 19 9 5 QMOD
Q2N 4 7 5 QMOD ;OFF
QSC 4 12 8 QMOD ;OFF
QOUT 19 1 11 QOUT 10
FEE 5 21 VCHAIN 6
EREF 6 21 15 21 5
FX 21 15 VCHAIN 1
VCHAIN 16 2 0
FAP 3 19 VCHAIN 300M
JON 2 21 21 JMOD
JST 19 21 21 JSTMOD
DBLK 21 19 DBLK ;OFF
DXX 19 16 DMOD
DREF 13 9 DMOD
DAP 3 19 DMOD ;OFF
DSC 12 14 DSCMOD ;OFF
DOUT 4 1 DMOD
RBLK 21 19 50K
RX 21 15 10K TC=0,-1040N
RSS 6 9 20
RDD 13 19 1MEG
ROMP 7 10 890
RZZ 8 7 5K
RSC2 14 19 40K
R2 21 8 5K
RAP 4 19 2MEG
RXX 12 11 530
RM 11 1 200K
RSC 8 11 0.27
CC2 7 21 0.7N
C_OMP 4 10 0.35N

.MODEL QMOD NPN IS=10F 
.MODEL QSCMOD NPN IS=10F NF=1.1 NR=1.1 
.MODEL JMOD NJF VTO=-4 BETA=6.25U 
.MODEL JSTMOD NJF VTO=-4 BETA=147.8125U 
.MODEL DMOD D 
.MODEL QPMOD PNP IS=10F BF=10 
.MODEL QOUT NPN IS=10F BF=10K RE=0.1 
.MODEL DBLK D BV=50 
.MODEL DSCMOD D BV=7 
.ENDS LM7805C

Rout OUT 0 1.0E3  
X1I6 IN OUT 0 LM7805C  
V1I41 IN 0 DC 10.0 AC 0.0  
.TRAN 0.1M 10M
.END

