RCL

R1 N2 N3 10.0  
L1 N2 N1 10.0E-3  
L2 N3 N4 10.0E-3  
V1I95 N1 0 AC 0.0 SIN ( 0.0 5.0 1.0E3 0.0 0.0 0.0 )  
R2 0 N4 10.0  
C1 N2 N4 10.0E-6  

.TRAN 0.1M 10M
.LIB
.IC V(2)=3 V(2)=4
.END

