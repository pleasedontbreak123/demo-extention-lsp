jfet_test
.MODEL N3972_LOW_SPEED NJF ( VTO=-1.12
+ BETA=10.6M LAMBDA=28.1M RD=4.37 RS=2.39 
+ CGS=23.4P CGD=23.4P PB=0.5 IS=1.846P )

V1 G1 0 AC 0.0 SIN ( 0.0 1.0 1.0E3 0.0 0.0 0.0 )  
V2 D1 0 AC 0.0 SIN ( 0.0 1.0 1.0E3 0.0 0.0 0.0 )  
RB G1 G 1.0E3  
RE S 0 1.0E3  
RC D1 D 10.0E3  
J1 D G S N3972_LOW_SPEED

.TRAN 1U 10M
.END