.SUBCKT one
R1 1 1 1

.SUBCKT two
R2 1 1 1
.ENDS two

.SUBCKT one
R3 1 1 1
.ENDS one

R4 1 1 1
.ENDS one
