
.option uselastdef

.MODEL 2N2222 NPN ( IS=39.4876F 
+ BF=200.9555 NF=1.0156 VAF=45.0913 IKF=2.9481 
+ ISE=0.1147P NE=1.4807 BR=18.0396 NR=1.0161 
+ VAR=10.0311 IKR=0.144 ISC=22.8562P NC=1.6619 
+ RB=5 IRB=54.3528U RBM=1.0644 RE=0.4936 
+ RC=0.6048 CJE=26.686P VJE=0.7111 MJE=0.332 
+ TF=0.1353N XTF=2 ITF=0.1576 CJC=14.2045P 
+ VJC=0.5142 MJC=0.3308 TR=16.5009N EG=1.11 )

.model a2d_eldo a2d mode=std_logic
.model d2a_eldo d2a mode=std_logic TRISE=50e-12 TFALL=50e-12
.defhook a2d_eldo
.defhook d2a_eldo
Q1I1 R2 N1N21 N1N260 2n2222  
R1 V1 N1N21 0.001  
C1 N1N21 0 1.0E-10  
V1 V1 0 AC 0.0 SIN ( 0.0 0.2 2.0E8 0.0 1.0E-9 0.0 )  
C2 R2 0 1.0E-10  
R2 N1N252 R2 100.0  
V2 N1N252 0 AC 0.0 PULSE ( 0.0 15.0 0.0 1.0E-9 1.0E-9 95.0 100.0 )  
C4 R4 0 1.0E-10  
Q1I146 R4 N1N257 N1N260 2n2222  
R3 N1N257 0 0.001  
C3 N1N257 0 1.0E-10  
C5 N1N260 0 1.0E-10  
R4 N1N252 R4 100.0  
I1I278 N1N260 0 AC 0.0 PULSE ( 0.0 0.16 0.0 1.0E-9 1.0E-9 95.0 100.0 )  
* Dictionary 1
* GND = 0
*.END
*Globals
