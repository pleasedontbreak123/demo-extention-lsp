R6

R1 1 2 1
R2 1 3 1
R3 5 4 1
R4 3 4 1
R5 2 3 1
R6 4 6 1
Vus1 1 6 DC 5
Vus2 2 5 DC 5

.control
  tran 0.1ms 10ms     
  plot v(1) v(2) v(4) v(5) v(6)    
.endc

.TRAN 1M 1 
.END
