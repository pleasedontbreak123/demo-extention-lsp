* Design ctr_sourse
* AMS Spice Netlist
* File created Mon Oct 14 15:24:31 2024
* ConfigFile:  C:\MentorGraphics\EEVX.2.8\SDD_HOME\standard\svspice.cfg
* Options   :  -60 -_ -h -kC:\MentorGraphics\EEVX.2.8\SDD_HOME\standard\svspice.cfg -gctr_sourse.tempfile ctr_sourse
*
.option uselastdef
* These libraries are listed in the [SpiceLibs] section
* of svnetlister.ini
*
*
* end of [SpiceLibs] section.
.MODEL 1N4001 D ( IS=11.4956P 
+ RS=0.114 N=1.321 CJO=36.1697P VJ=0.583 
+ M=0.464 BV=50 IBV=50N )

.model a2d_eldo a2d mode=std_logic
.model d2a_eldo d2a mode=std_logic TRISE=50e-12 TFALL=50e-12
.defhook a2d_eldo
.defhook d2a_eldo
V1I251 VIN 0 DC 5.0 AC 0.0 0.0  
V1I175 VCTR 0 AC 0.0 SIN ( 1.0 1.0 1.0E3 0.0 0.0 0.0 )  
E1I242 VIN VOUT VCTR 0 1.0  
G1I266 IIN IOUT VCTR 0 1.0  
R1I176 VOUT 0 1.0E3  
R1I313 VIN IIN 1.0E3  
Dd1 0 IOUT 1N4001  
H1I321 VIN VOUT2 Vsin 1.0  
Vsin ICTR 0 AC 0.0 SIN ( 0.0 1.0 1.0E3 0.0 0.0 0.0 )  
R1I347 VOUT2 0 1.0E3  
Rr1 0 ICTR 1.0E3  
F1I452 IIN2 IOUT2 Vsin 1.0  
Rout IOUT2 0 1.0E3  
I1I506 IIN2 N1N492 DC 5.0 AC 1.0  
R1I493 IIN2 N1N492 1.0E3  
* Dictionary 10
* Iout2=IOUT2
* Iin2=IIN2
* Ictr=ICTR
* Vout2=VOUT2
* Iout=IOUT
* Iin=IIN
* Vout=VOUT
* Vctr=VCTR
* GND=0
* Vin = VIN
*.END
*Globals
