* Design figure5
* AMS Spice Netlist
* File created Mon Sep 30 10:32:43 2024
* ConfigFile:  C:\MentorGraphics\EEVX.2.8\SDD_HOME\standard\svspice.cfg
* Options   :  -60 -_ -h -kC:\MentorGraphics\EEVX.2.8\SDD_HOME\standard\svspice.cfg -gfigure5.tempfile figure5
*
.option uselastdef
* These libraries are listed in the [SpiceLibs] section
* of svnetlister.ini
*
*
* end of [SpiceLibs] section.
.MODEL DSK10C          D ( IS=2.729e-07 
+ RS=0.0298 N=2.422 TT=1e-10 CJO=1e-13 
+ VJ=1 BV=200 IBV=0.001 EG=1.11 
+ XTI=5 KF=0 AF=1 FC=0.5 
+ M=0.5 )
.subckt vc_sw_spice np nn cp cn PARAM: level=1 von=0.95 voff=0.05 ron=0.05 roff=100.0e3
YSW vswitch np nn cp cn PARAM: level=level von=von voff=voff ron=ron roff=roff MODEL: vc_sw
.model vc_sw modfas
.ends
* Models for Eldo<->VHDL-AMS data conversion
.model a2d_eldo a2d mode=std_logic
.model d2a_eldo d2a mode=std_logic TRISE=50e-12 TFALL=50e-12
.defhook a2d_eldo
.defhook d2a_eldo
V1I239 IN 0 DC 24.0 AC 0.0  
V1I263 N1N296 0 AC 0.0 PULSE ( 0.0 1.0 0.0 0.01E-3 0.01E-3 0.1E-3 0.2E-3 )  
Ll1 N1 OUT 0.1E-3  
C1I69 OUT 0 0.1E-3  
R1I29 OUT 0 10.0  
D1I39 0 OUT DSK10C  
X1I257 IN N1 N1N296 0 vc_sw_spice LEVEL=1.0 ROFF=100000.0 RON=0.00001 VOFF=0.05 
+ VON=0.5  
* Dictionary 4
* out=OUT
* 1=N1
* GND=0
* in = IN
*.END
*Globals
